module example (
// Clock and active low Asynchronous Reset
    input logic clk,rst_n 
// Signals    
    //,
);
// Enter your code here
endmodule
